//`define REG_PROTECTION_HAMMING
`define REG_PROTECTION_HAMMING
`define USE_UNPROTECTED_PART
