`define REG_PROTECTION_MJR
`define USE_UNPROTECTED_PART