/*
`ifndef CRC_MACRO

`define CRC_MACRO

//`define REG_PROTECTION_HAMMING
`define REG_PROTECTION_MJR

`endif //CRC_MACRO*/
