`define REG_PROTECTION_MJR
`define FORCE_MJR_REG
`define FORCE_REGISTER_PROTECTION
