
`ifndef CRC_MACRO

`define CRC_MACRO

`define REG_PROTECTION_HAMMING

`endif //CRC_MACRO
